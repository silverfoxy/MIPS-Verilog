library verilog;
use verilog.vl_types.all;
entity Core_TB is
end Core_TB;
